
module test();


    woof
     





    
    
endmodule 
