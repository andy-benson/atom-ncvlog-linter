
module test();


    woof
     







    
    
endmodule 
