module lint_test();
   


   wire woof;
   wire jjdjjd


   assign woof             = 1'b1;
   assign woofjdhjsahdjahdjkakd = 1'b1;


endmodule 
